//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// SystemVerilog version Alex Grinshpun May 2018
// coding convention dudy December 2018
// (c) Technion IIT, Department of Electrical Engineering 2019 


module	back_ground_drawSquare	(	

					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0]	pixelX,
					input logic	[10:0]	pixelY,
					input logic startOfFrame,
					input logic pause,
					output	logic	[7:0]	BG_RGB
);

parameter int BG_SPEED = 148;

logic [0:31] offsetFIXED;

logic [0:5] offset;

const int FIXED_POINT_MULIPLIER=64;

localparam  int OBJECT_HEIGHT_Y = 64;
localparam  int OBJECT_WIDTH_X = 64;

logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors = {
{8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75 },
{8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75 },
{8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'h99, 8'h99, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51 },
{8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'h99, 8'h99, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51 },
{8'h99, 8'h99, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51 },
{8'h99, 8'h99, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51 },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51 },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51 },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD },
{8'hBD, 8'hBD, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'hBD, 8'hBD, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'hBD, 8'hBD, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'hBD, 8'hBD, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'hBD, 8'hBD, 8'h75, 8'h75, 8'h99, 8'h99, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h99, 8'h99, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'hBD, 8'hBD, 8'h75, 8'h75, 8'h99, 8'h99, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h99, 8'h99, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD },
{8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD },
{8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h99, 8'h99, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD },
{8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h99, 8'h99, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD },
{8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h51, 8'h51, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'hBD, 8'hBD, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h51, 8'h51, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'hBD, 8'hBD, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h99, 8'h99, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h99, 8'h99, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51 },
{8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51 },
{8'h75, 8'h75, 8'h51, 8'h51, 8'h99, 8'h99, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51 },
{8'h75, 8'h75, 8'h51, 8'h51, 8'h99, 8'h99, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51 },
{8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51 },
{8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51 },
{8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51 },
{8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51 },
{8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h50, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h51, 8'h51 },
{8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h50, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h51, 8'h51 },
{8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'hBD, 8'hBD, 8'h51, 8'h51 },
{8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'h51, 8'h51, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'hBD, 8'hBD, 8'h51, 8'h51 },
{8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'h50, 8'h50, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75 },
{8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h30, 8'h30, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h30, 8'h30, 8'h50, 8'h50, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD },
{8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD },
{8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h99, 8'h99 },
{8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h99, 8'h99 },
{8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h50, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99 },
{8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h50, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99 },
{8'h50, 8'h50, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h50, 8'h50, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h50, 8'h50, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h50, 8'h50, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h99, 8'h99, 8'h51, 8'h51, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75 },
{8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50 },
{8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h50, 8'h50 },
{8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C },
{8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h51, 8'h51, 8'h50, 8'h50, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h30, 8'h30, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h2C, 8'h2C },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C },
{8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h75, 8'h2C, 8'h2C, 8'h51, 8'h51, 8'h75, 8'h75, 8'h99, 8'h99, 8'h51, 8'h51, 8'h2C, 8'h2C, 8'hBD, 8'hBD, 8'h75, 8'h75, 8'h50, 8'h50, 8'h51, 8'h51, 8'h75, 8'h75, 8'h75, 8'h75, 8'h99, 8'h99, 8'h75, 8'h75, 8'h2C, 8'h2C }
};


const int	xFrameSize	=	639;
const int	yFrameSize	=	479;

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		BG_RGB <= object_colors[pixelY][pixelX];
	end 
	else begin	

		if(pause) 	begin
			BG_RGB <= object_colors[pixelY-offset][pixelX];
			offsetFIXED<=offsetFIXED;
		end
		else begin
			BG_RGB <= object_colors[pixelY-offset][pixelX];
			if (startOfFrame) offsetFIXED<=offsetFIXED+BG_SPEED;
		end
	
	end; 	
end

assign offset = offsetFIXED/FIXED_POINT_MULIPLIER;
 
endmodule

