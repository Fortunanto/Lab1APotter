////-- Alex Grinshpun Apr 2017
////-- Dudy Nov 13 2017
//// System-Verilog Alex Grinshpun May 2018
//// New coding convention dudy December 2018
//// (c) Technion IIT, Department of Electrical Engineering 2019 
//
//
//module	towers_moveCollision	(	
//					input		logic	clk,
//					input		logic	resetN,
//					input    logic startOfFrame,
//					
//					input shortint score,
//					
//					//output   logic edgeCollide,
//					output	logic	drawingRequest // indicates pixel inside the bracket				
//);
//
//parameter int DIGITS_AMOUNT = 5;
//
//logic [0:DIGITS_AMOUNT-1][0:3] digits;
//
//genvar i;
//generate
//	for (i=0;i<DIGITS_AMOUNT;i++) begin: digigen
//		
//	end
//endgenerate
//
//endmodule 