module shot_soundModulator();
endmodule